library verilog;
use verilog.vl_types.all;
entity t_1017_3 is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        W               : out    vl_logic_vector(5 downto 0)
    );
end t_1017_3;
