`timescale 1ns/10ps
module counter_4bit_0_5(
	input reset,					//重置
	input clk,						//時脈
	input carry_in, 				//進位輸入
	output logic [3:0] value, 	//輸出
	output logic carry_out 		//進位輸出
);

	always_ff @ (posedge clk)
		begin
			if(reset)              //同步，如果reset 就把值歸0
				value <= #1 0;
			else if(value == 4'd5 && carry_in == 1) //數到5也把值歸0
				value <= #1 0;
			else if(carry_in == 1)
				value <= #1 value + 1; //值加1
		end
		
	assign carry_out = (value == 4'd5 && carry_in == 1)?1:0; //當value = 5 且 carry_in = 1時，有進位
	
endmodule